
module x;



parameter AA = 2;

if (AA>2) begin
    wire [3:0] [5:0] xxx;
end


endmodule

